`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    15:00:38 11/23/2016 
// Design Name: 
// Module Name:    ControllerM 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module ControllerM(
    input [5:0] Op,
    output MemWrite
    );
	assign MemWrite = Op == 101011; //sw

endmodule
